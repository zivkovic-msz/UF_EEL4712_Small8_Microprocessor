library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity internal_architecture is
	generic ( 
		width : positive := 8);
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end internal_architecture;

architecture STR of internal_architecture is







end STR;