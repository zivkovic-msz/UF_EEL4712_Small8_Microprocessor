library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity alu_tb is
end alu_tb;

architecture TB of alu_tb is

    constant WIDTH  : positive := 8;
	signal input_A	: std_logic_vector(WIDTH-1 downto 0) := (others => '0');
	signal input_D	: std_logic_vector(WIDTH-1 downto 0) := (others => '0');
	signal sel		: std_logic_vector(3 downto 0) := (others => '0');
	signal output	: std_logic_vector(WIDTH-1 downto 0) := (others => '0');
	signal carry_in : std_logic_vector(0 downto 0) := (others => '0');
	signal carry_flag : std_logic_vector(0 downto 0) := (others => '0');
	signal overflow_flag : std_logic_vector(0 downto 0) := (others => '0'); 
	signal signed_flag : std_logic_vector(0 downto 0) := (others => '0');
	signal zero_flag : std_logic_vector(0 downto 0) := (others => '0');

begin  -- TB

    UUT : entity work.alu
        generic map (WIDTH => WIDTH)
        port map (
            input_A  => input_A,
            input_D   => input_D,
            sel      => sel,
            output   => output,
			carry_in => carry_in,
			carry_flag => carry_flag,
			overflow_flag => overflow_flag,
			signed_flag => signed_flag,
			zero_flag => zero_flag 
            );

    process
    begin
		
		--Test zero flag
		sel    <= "0000";
		carry_in(0) <= '0';
        input_A <= conv_std_logic_vector(0, input_A'length);
        input_D <= conv_std_logic_vector(0, input_D'length);
        wait for 40 ns;
		
        -- Add with carry overflow
        sel    <= "0000";
		carry_in(0) <= '1';
        input_A <= conv_std_logic_vector(250, input_A'length);
        input_D <= conv_std_logic_vector(50, input_D'length);
        wait for 40 ns;
		
        -- Add with carry overflow
        sel    <= "0000";
		carry_in(0) <= '1';
        input_A <= conv_std_logic_vector(250, input_A'length);
        input_D <= conv_std_logic_vector(5, input_D'length);
        wait for 40 ns;
		
		-- Add with carry no overflow
		sel    <= "0000";
		carry_in(0) <= '1';
       input_A <= conv_std_logic_vector(250, input_A'length);
       input_D <= conv_std_logic_vector(2, input_D'length);
       wait for 40 ns;
       
		--Subtract with borrow (overflow) (-112 - 96) = (1) 00110000 = 48
 		sel    <= "0001";
		carry_in(0) <= '1';
       input_A <= conv_std_logic_vector(-112, input_A'length); 
       input_D <= conv_std_logic_vector(96, input_D'length);
       wait for 40 ns;

		--Subtract with borrow (no overflow)
 		sel    <= "0001";
		carry_in(0) <= '1';
       input_A <= conv_std_logic_vector(7, input_A'length); 
       input_D <= conv_std_logic_vector(3, input_D'length);
       wait for 40 ns;
		
		-- Compare
		sel    <= "0010";
		carry_in(0) <= '1';
       input_A <= conv_std_logic_vector(5, input_A'length);
       input_D <= conv_std_logic_vector(4, input_D'length);
       wait for 40 ns;
		
		-- Compare
		sel    <= "0010";
		carry_in(0) <= '1';
       input_A <= conv_std_logic_vector(5, input_A'length);
       input_D <= conv_std_logic_vector(5, input_D'length);
       wait for 40 ns;
		
		--AND
		sel    <= "0011";
		carry_in(0) <= '1';
        input_A <= conv_std_logic_vector(255, input_A'length);
        input_D <= conv_std_logic_vector(170, input_D'length);
        wait for 40 ns;
		
		--OR
		sel    <= "0100";
		carry_in(0) <= '1';
        input_A <= conv_std_logic_vector(255, input_A'length);
        input_D <= conv_std_logic_vector(170, input_D'length);
        wait for 40 ns;
		
		--XOR
		sel    <= "0101";
		carry_in(0) <= '1';
        input_A <= conv_std_logic_vector(255, input_A'length);
        input_D <= conv_std_logic_vector(170, input_D'length);
        wait for 40 ns;
		
		--Shift Left Logical
		sel    <= "0110";
        input_A <= conv_std_logic_vector(212, input_A'length);
        input_D <= conv_std_logic_vector(0, input_D'length);
        wait for 40 ns;		
		
		--Shift Right Logical
		sel    <= "0111";
        input_A <= conv_std_logic_vector(212, input_A'length);
        input_D <= conv_std_logic_vector(0, input_D'length);
        wait for 40 ns;		
		
		--Rotate Left through Carry
		sel    <= "1000";
		carry_in(0) <= '1';
        input_A <= conv_std_logic_vector(212, input_A'length);
        input_D <= conv_std_logic_vector(0, input_D'length);
        wait for 40 ns;		
		
		--Rotate Right through Carry
		sel    <= "1001";
		carry_in(0) <= '1';
        input_A <= conv_std_logic_vector(212, input_A'length);
        input_D <= conv_std_logic_vector(0, input_D'length);
        wait for 40 ns;			
		
		--Decrement Acc
		sel    <= "1010";
        input_A <= conv_std_logic_vector(15, input_A'length);
        input_D <= conv_std_logic_vector(0, input_D'length);
        wait for 40 ns;		
		
		--Increment Acc
		sel    <= "1011";
        input_A <= conv_std_logic_vector(15, input_A'length);
        input_D <= conv_std_logic_vector(0, input_D'length);
        wait for 40 ns;
		
		--Set Carry Flag
		sel    <= "1100";
        wait for 40 ns;		
		
		--Clear Carry Flag
		sel    <= "1101";
        wait for 40 ns;				
		
		
        -- test 250+50 (with overflow)
		-- -- carry_in <= '
        -- -- sel    <= "0000";
        -- -- input_A <= conv_std_logic_vector(250, input_A'length);
        -- -- input_D <= conv_std_logic_vector(50, input_D'length);
        -- -- wait for 40 ns;
       -- assert(output = conv_std_logic_vector(300, output'length)) report "Error : 250+50 = " & integer'image(conv_integer(output)) & " instead of 44" severity warning;
       -- assert(overflow = '1') report "Error                                     : overflow incorrect for 250+50" severity warning;


		-- test subtraction
		-- -- sel    <= "0001";
		-- -- carry_in <= '1';
        -- -- input_A <= conv_std_logic_vector(15, input_A'length);
        -- -- input_D <= conv_std_logic_vector(10, input_D'length);
        -- -- wait for 40 ns;
       -- assert(output = conv_std_logic_vector(5, output'length)) report "Error : 15-10 = " & integer'image(conv_integer(output)) & " instead of 5" severity warning;
       -- assert(overflow = '0') report "Error overflow incorrect." severity warning;

		
        -- test 5*6
        -- -- sel    <= "0010";
        -- -- input_A <= conv_std_logic_vector(5, input_A'length);
        -- -- input_D <= conv_std_logic_vector(6, input_D'length);
        -- -- wait for 40 ns;
        -- -- assert(output = conv_std_logic_vector(30, output'length)) report "Error : 5*6 = " & integer'image(conv_integer(output)) & " instead of 30" severity warning;
        -- -- assert(overflow = '0') report "Error                                    : overflow incorrect for 5*6" severity warning;

        -- test 50*60
        -- -- sel    <= "0010";
        -- -- input_A <= conv_std_logic_vector(64, input_A'length);
        -- -- input_D <= conv_std_logic_vector(64, input_D'length);
        -- -- wait for 40 ns;
        -- -- assert(output = conv_std_logic_vector(4096, output'length)) report "Error : 64*64 = " & integer'image(conv_integer(output)) & " instead of 0" severity warning;
        -- -- assert(overflow = '1') report "Error                                      : overflow incorrect for 64*64" severity warning;

        -- test AND
        -- -- sel <= "0011";
        -- -- input_A <= conv_std_logic_vector(15, input_A'length);
        -- -- input_D <= conv_std_logic_vector(10, input_D'length);
        -- -- wait for 40 ns;
        -- -- assert(output = conv_std_logic_vector(10, output'length)) report "Error : 0xF AND 0xA = " & integer'image(conv_integer(output)) & " instead of 0xA" severity warning;
        -- -- assert(overflow = '0') report "Error                                    : overflow incorrect for 0xF AND 0xA" severity warning;  
        
        -- test OR
        -- -- sel <= "0100";
        -- -- input_A <= conv_std_logic_vector(15, input_A'length);
        -- -- input_D <= conv_std_logic_vector(10, input_D'length);
        -- -- wait for 40 ns;
        -- -- assert(output = conv_std_logic_vector(15, output'length)) report "Error : 0xF OR 0xA = " & integer'image(conv_integer(output)) & " instead of 0xF" severity warning;
        -- -- assert(overflow = '0') report "Error : overflow incorrect" severity warning;
        
        -- test XOR
        -- -- sel <= "0101";
        -- -- input_A <= conv_std_logic_vector(15, input_A'length);
        -- -- input_D <= conv_std_logic_vector(10, input_D'length);
        -- -- wait for 40 ns;
        -- -- assert(output = conv_std_logic_vector(5, output'length)) report "Error : 0xF XOR 0xA = " & integer'image(conv_integer(output)) & " instead of 0x5" severity warning;
        -- -- assert(overflow = '0') report "Error : overflow incorrect" severity warning;
        
        -- test NOR
        -- -- sel <= "0110";
        -- -- input_A <= conv_std_logic_vector(15, input_A'length);
        -- -- input_D <= conv_std_logic_vector(10, input_D'length);
        -- -- wait for 40 ns;
        -- -- assert(output(3 downto 0) = "0000") report "Error : 0xF NOR 0xA = " & integer'image(conv_integer(output)) & " instead of 0x0" severity warning;
        -- -- assert(overflow = '0') report "Error : overflow incorrect" severity warning;
        
        -- test NOT
        -- -- sel <= "0111";
        -- -- input_A <= conv_std_logic_vector(9, input_A'length);
        -- input_D <= conv_std_logic_vector("1010", input_D'length);
        -- -- wait for 40 ns;
        -- -- assert(output(3 downto 0) = "0110") report "Error : NOT 0x9 = " & integer'image(conv_integer(output)) & " instead of 0x6" severity warning;
        -- -- assert(overflow = '0') report "Error : overflow incorrect" severity warning;
        
        -- test Shift left 1 bit
        -- -- sel <= "1000";
        -- -- input_A <= conv_std_logic_vector(11, input_A'length);
        -- input_D <= conv_std_logic_vector("1010", input_D'length);
        -- -- wait for 40 ns;
       -- assert(output = conv_std_logic_vector(6, output'length)) report "Error : SHIFT_LEFT(1011) = " & integer'image(conv_integer(output)) & " instead of 0110" severity warning;
        -- -- if(input_A(WIDTH-1) = '1') then
        -- -- assert(overflow = '1') report "Error : overflow incorrect" severity warning;
        -- -- end if;
        
        -- test shift right 1 bit
        -- -- sel <= "1001";
        -- -- input_A <= conv_std_logic_vector(11, input_A'length); --1011
        -- input_D <= conv_std_logic_vector("1010", input_D'length);
        -- -- wait for 40 ns;
        -- -- assert(output = conv_std_logic_vector(5, output'length)) report "Error : SHIFT_RIGHT(1011) = " & integer'image(conv_integer(output)) & " instead of 0101" severity warning;
        -- -- assert(overflow = '0') report "Error : overflow incorrect" severity warning;             
        
        -- test swap
        -- -- sel <= "1010";
        -- -- input_A <= conv_std_logic_vector(40, input_A'length); --101000
        -- input_D <= conv_std_logic_vector("1010", input_D'length);
        -- -- wait for 40 ns;
        -- assert(output = conv_std_logic_vector(5, output'length)) report "Error : swap = " & integer'image(conv_integer(output)) & " instead of 0000101" severity warning;
        -- -- assert(overflow = '0') report "Error : overflow incorrect" severity warning;    

        -- test reverse bits
        -- -- sel <= "1011";
        -- -- input_A <= conv_std_logic_vector(10, input_A'length);
        -- input_D <= conv_std_logic_vector("1010", input_D'length);
        -- -- wait for 40 ns;
        -- assert(output = conv_std_logic_vector(5, output'length)) report "Error : reverse bits = " & integer'image(conv_integer(output)) & " instead of 0101" severity warning;
        -- -- assert(overflow = '0') report "Error : overflow incorrect" severity warning;  
        
        -- test other select bits
        -- -- sel <= "1100";
        -- -- input_A <= "01101011";
        -- -- wait for 40 ns;
        -- assert(output = conv_std_logic_vector(0,output'length)) report "Error, output should  be 0" severity warning;
        -- -- sel <= "1101";
        -- -- input_D <= "00000011";
        -- -- input_A <= "00000010";
        -- -- wait for 40 ns;
        -- assert(output = conv_std_logic_vector(0,output'length)) report "Error, output should  be 0" severity warning;
        -- -- sel <= "1110";
        -- -- input_A <= "10101010";
        -- -- input_D <= "10101010";
        -- -- wait for 40 ns;
        -- assert(output = conv_std_logic_vector(0,output'length)) report "Error, output should  be 0" severity warning;
        -- -- sel <= "1111";
        -- -- input_A <= "01101011";
        -- -- wait for 40 ns;
        -- assert(output = conv_std_logic_vector(0,output'length)) report "Error, output should  be 0" severity warning;
        
        wait;

    end process;

end TB;
